library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use IEEE.NUMERIC_STD.ALL;
use IEEE.MATH_REAL.ALL;

Entity SRA64 is
Generic ( N : natural := 64 );
Port ( X : in std_logic_vector( N-1 downto 0 );
	Y : out std_logic_vector( N-1 downto 0 );
	ShiftCount : in unsigned( integer(ceil(log2(real(N))))-1 downto 0 ) );
End Entity SRA64;

Architecture rtl of SRA64 is 
	signal Y1, Y2, Y3 : std_logic_vector(N-1 downto 0);
	signal signExt: std_logic_vector(N-1 downto 0);
	signal shiftCountBits: std_logic_vector(5 downto 0);
Begin
	shiftCountBits <= std_logic_vector(ShiftCount);
	
	--First Barrel Shifter for SRA of 0, 16, 32, 48
	Y1 <= 	x"0000" & X(N-1 downto 16) when shiftCountBits(5 downto 4) = "01" else 
		x"00000000" & X(N-1 downto 32) when shiftCountBits(5 downto 4) = "10" else 
		x"000000000000" & X(N-1 downto 48) when shiftCountBits(5 downto 4) = "11" else 
		X;

	--Second Barrel Shifter for SRA of 0, 4, 8, 12
	Y2 <= 	x"0" & Y1(N-1 downto 4) when shiftCountBits(3 downto 2) = "01" else 
		x"00" & Y1(N-1 downto 8)  when shiftCountBits(3 downto 2) = "10" else 
		x"000" & Y1(N-1 downto 12) when shiftCountBits(3 downto 2) = "11" else 
		Y1;

	--Third Barrel Shifter for SRA of 0, 1, 2, 3
	Y3 <= 	"0" & Y2(N-1 downto 1) when shiftCountBits(1 downto 0) = "01" else 
		"00" & Y2(N-1 downto 2) when shiftCountBits(1 downto 0) = "10" else 
		"000" & Y2(N-1 downto 3) when shiftCountBits(1 downto 0) = "11" else 
		Y2;

	signExt(N-1-to_integer(ShiftCount) downto 0) <= Y3(N-1-to_integer(ShiftCount) downto 0); 
	signExt(N-1 downto N-to_integer(ShiftCount)) <= (N-1 downto N-to_integer(ShiftCount) => Y3(N-to_integer(ShiftCount)));
	Y <= signExt;

End Architecture rtl;